module Register_IF_ID
(
    instr_i,
    instrAddr_i,
    IFIDWrite_i,
    IFFlush_i,
    instr_o,
    instrAddr_o
);

// Interface


// Calculate

endmodule
