module Hazard_Detection_Unit
(
    ID_rsAddr_i,
    ID_rtAddr_I,
    EX_memRead_i,
    EX_wbAddr_i,
    hazardDetected_i
);

// Interface

// Calculation


endmodule