module WB_Addr_MUX
(
    rtAddr_i,
    rdAddr_i,
    wbDst_i,
    wbAddr_o
);

// Interface

// Calculation


endmodule
