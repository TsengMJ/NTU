module Sign_Extend
(
    imm_i,
    immExtended_o
);


// Interface


// Calculate

endmodule
