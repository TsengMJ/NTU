`define CYCLE_TIME 50            
`include "CPU.v"

module TestBench;

reg                Clk;
reg                Start;
integer            i, outfile, counter;
integer            stall, flush;

always #(`CYCLE_TIME/2) Clk = ~Clk;    


CPU CPU(
    .clk_i  (Clk),
    .start_i(Start)
);
  
initial begin
    $dumpfile("Project_1.vcd");
    $dumpvars;
    
    counter = 0;
    stall = 0;
    flush = 0;
    
    // initialize instruction memory
    for(i=0; i<256; i=i+1) begin
        CPU.Instruction_Memory.memory[i] = 32'b0;
    end
    
    // initialize data memory
    for(i=0; i<32; i=i+1) begin
        CPU.Data_Memory.memory[i] = 8'b0;
    end    

    // initialize Register File
    for(i=0; i<32; i=i+1) begin
        CPU.Registers.register[i] = 32'b0;
    end

    // initialize PC register
    CPU.PC.pc_o = 32'b0;

    // TODO: initialize pipeline registers
<<<<<<< HEAD:Classes/Computer_Architecture/HW/4/code/testbench.v
    	CPU.Register_IF_ID.instr_o = 32'b0;
	CPU.Register_IF_ID.instrAddr_o = 32'b0;

	CPU.Register_ID_EX.rsData_o= 32'b0;
	CPU.Register_ID_EX.rtData_o= 32'b0;
	CPU.Register_ID_EX.immExtended_o= 32'b0;
	CPU.Register_ID_EX.aluOp_o= 2'b0;
	CPU.Register_ID_EX.aluSrc_o= 1'b0;
	CPU.Register_ID_EX.wbDst_o= 1'b0;
	CPU.Register_ID_EX.memRead_o= 1'b0;
	CPU.Register_ID_EX.memWrite_o= 1'b0;
	CPU.Register_ID_EX.memToReg_o= 1'b0;
	CPU.Register_ID_EX.regWrite_o= 1'b0;
	CPU.Register_ID_EX.rsAddr_o= 4'b0;
	CPU.Register_ID_EX.rtAddr_o= 4'b0;
	CPU.Register_ID_EX.rdAddr_o= 4'b0;
	CPU.Register_ID_EX.funct_o= 10'b0;


	CPU.Register_EX_MEM.aluResult_o= 32'b0;
	CPU.Register_EX_MEM.aluSrc2_o	= 32'b0;
	CPU.Register_EX_MEM.memRead_o= 1'b0;
	CPU.Register_EX_MEM.memWrite_o= 1'b0;
	CPU.Register_EX_MEM.memToReg_o= 1'b0;
	CPU.Register_EX_MEM.regWrite_o= 1'b0;
	CPU.Register_EX_MEM.wbAddr_o= 6'b0;

	CPU.Register_MEM_WB.memData_o= 32'b0;
	CPU.Register_MEM_WB.aluResult_o= 32'b0;
	CPU.Register_MEM_WB.memToReg_o= 1'b0;
	CPU.Register_MEM_WB.regWrite_o= 1'b0;
	CPU.Register_MEM_WB.wbAddr_o  = 6'b0;
=======
    CPU.Hazard_Detection_Unit.hazardDetected_o = 1'b0;
    CPU.Register_IF_ID.instr_o = 32'b0;
	CPU.Register_IF_ID.instrAddr_o = 32'b0;

	CPU.Register_ID_EX.rsData_o = 32'b0;
	CPU.Register_ID_EX.rtData_o = 32'b0;
	CPU.Register_ID_EX.immExtended_o = 32'b0;
	CPU.Register_ID_EX.aluOp_o = 2'b0;
	CPU.Register_ID_EX.aluSrc_o = 1'b0;
	CPU.Register_ID_EX.memRead_o = 1'b0;
	CPU.Register_ID_EX.memWrite_o = 1'b0;
	CPU.Register_ID_EX.memToReg_o = 1'b0;
	CPU.Register_ID_EX.regWrite_o = 1'b0;
	CPU.Register_ID_EX.rsAddr_o = 5'b0;
	CPU.Register_ID_EX.rtAddr_o = 5'b0;
	CPU.Register_ID_EX.rdAddr_o = 5'b0;
    CPU.Register_ID_EX.wbAddr_o = 5'b0;
	CPU.Register_ID_EX.funct_o = 10'b0;


    

	CPU.Register_EX_MEM.aluResult_o = 32'b0;
	CPU.Register_EX_MEM.rtData_o = 32'b0;
	CPU.Register_EX_MEM.memRead_o = 1'b0;
	CPU.Register_EX_MEM.memWrite_o = 1'b0;
	CPU.Register_EX_MEM.memToReg_o = 1'b0;
	CPU.Register_EX_MEM.regWrite_o = 1'b0;
	CPU.Register_EX_MEM.wbAddr_o = 5'b0;

	CPU.Register_MEM_WB.memData_o = 32'b0;
	CPU.Register_MEM_WB.aluResult_o = 32'b0;
	CPU.Register_MEM_WB.memToReg_o = 1'b0;
	CPU.Register_MEM_WB.regWrite_o = 1'b0;
	CPU.Register_MEM_WB.wbAddr_o  = 5'b0;



    
>>>>>>> da8f5dc6281b5542f4b7345dab5f5a7e2bd8ab44:Classes/Computer_Architecture/HW/4/code (Ori)/testbench.v

    // Load instructions into instruction memory

    // $readmemb("../testdata/instruction.txt", CPU.Instruction_Memory.memory);
    $readmemb("../testdata/Fibonacci_instruction.txt", CPU.Instruction_Memory.memory);
    
    // Open output file
    outfile = $fopen("../testdata/output.txt") | 1;
    
    // Set Input n into data memory at 0x00
    CPU.Data_Memory.memory[0] = 8'h5;       // n = 5 for example
    
    Clk = 1;
    //Reset = 0;
    Start = 0;
    
    #(`CYCLE_TIME/4) 
    //Reset = 1;
    Start = 1;
        
    
end
  
always@(posedge Clk) begin
    // TODO: change # of cycles as you need
    // if(counter == 30)    // stop after 30 cycles
    //     $finish;
    if(counter == 64)    // stop after 30 cycles
        $finish;

    // TODO: put in your own signal to count stall and flush
    if(CPU.Hazard_Detection_Unit.hazardDetected_o == 1 && CPU.Control.branch_o == 0) stall = stall + 1;
    if(CPU.Control.flush_o == 1) flush = flush + 1;  
   

    // print PC
    $fdisplay(outfile, "cycle = %d, Start = %d, Stall = %d, Flush = %d\nPC = %d", counter, Start, stall, flush, CPU.PC.pc_o);
    
    // print Registers
    $fdisplay(outfile, "Registers");
    $fdisplay(outfile, "x0 = %d, x8  = %d, x16 = %d, x24 = %d", CPU.Registers.register[0], CPU.Registers.register[8] , CPU.Registers.register[16], CPU.Registers.register[24]);
    $fdisplay(outfile, "x1 = %d, x9  = %d, x17 = %d, x25 = %d", CPU.Registers.register[1], CPU.Registers.register[9] , CPU.Registers.register[17], CPU.Registers.register[25]);
    $fdisplay(outfile, "x2 = %d, x10 = %d, x18 = %d, x26 = %d", CPU.Registers.register[2], CPU.Registers.register[10], CPU.Registers.register[18], CPU.Registers.register[26]);
    $fdisplay(outfile, "x3 = %d, x11 = %d, x19 = %d, x27 = %d", CPU.Registers.register[3], CPU.Registers.register[11], CPU.Registers.register[19], CPU.Registers.register[27]);
    $fdisplay(outfile, "x4 = %d, x12 = %d, x20 = %d, x28 = %d", CPU.Registers.register[4], CPU.Registers.register[12], CPU.Registers.register[20], CPU.Registers.register[28]);
    $fdisplay(outfile, "x5 = %d, x13 = %d, x21 = %d, x29 = %d", CPU.Registers.register[5], CPU.Registers.register[13], CPU.Registers.register[21], CPU.Registers.register[29]);
    $fdisplay(outfile, "x6 = %d, x14 = %d, x22 = %d, x30 = %d", CPU.Registers.register[6], CPU.Registers.register[14], CPU.Registers.register[22], CPU.Registers.register[30]);
    $fdisplay(outfile, "x7 = %d, x15 = %d, x23 = %d, x31 = %d", CPU.Registers.register[7], CPU.Registers.register[15], CPU.Registers.register[23], CPU.Registers.register[31]);

    // print Data Memory
    $fdisplay(outfile, "Data Memory: 0x00 = %10d", {CPU.Data_Memory.memory[3] , CPU.Data_Memory.memory[2] , CPU.Data_Memory.memory[1] , CPU.Data_Memory.memory[0] });
    $fdisplay(outfile, "Data Memory: 0x04 = %10d", {CPU.Data_Memory.memory[7] , CPU.Data_Memory.memory[6] , CPU.Data_Memory.memory[5] , CPU.Data_Memory.memory[4] });
    $fdisplay(outfile, "Data Memory: 0x08 = %10d", {CPU.Data_Memory.memory[11], CPU.Data_Memory.memory[10], CPU.Data_Memory.memory[9] , CPU.Data_Memory.memory[8] });
    $fdisplay(outfile, "Data Memory: 0x0c = %10d", {CPU.Data_Memory.memory[15], CPU.Data_Memory.memory[14], CPU.Data_Memory.memory[13], CPU.Data_Memory.memory[12]});
    $fdisplay(outfile, "Data Memory: 0x10 = %10d", {CPU.Data_Memory.memory[19], CPU.Data_Memory.memory[18], CPU.Data_Memory.memory[17], CPU.Data_Memory.memory[16]});
    $fdisplay(outfile, "Data Memory: 0x14 = %10d", {CPU.Data_Memory.memory[23], CPU.Data_Memory.memory[22], CPU.Data_Memory.memory[21], CPU.Data_Memory.memory[20]});
    $fdisplay(outfile, "Data Memory: 0x18 = %10d", {CPU.Data_Memory.memory[27], CPU.Data_Memory.memory[26], CPU.Data_Memory.memory[25], CPU.Data_Memory.memory[24]});
    $fdisplay(outfile, "Data Memory: 0x1c = %10d", {CPU.Data_Memory.memory[31], CPU.Data_Memory.memory[30], CPU.Data_Memory.memory[29], CPU.Data_Memory.memory[28]});
	
    $fdisplay(outfile, "\n");
    
    counter = counter + 1;
    
      
end

  
endmodule
