module Register_EX_MEM
(
    memRead_i,
    memWrite_i,
    memToReg_i,
    aluResult_i,
    aluSrc2_i,
    wbAddr_i,

    memRead_o,
    memWrite_o,
    memToReg_o,
    aluResult_o,
    aluSrc2_o,
    wbAddr_o
);

// Interface

// Calculation


endmodule