module RT_IMM_MUX
(
    rtData_i,
    immExtended_i,
    alu_rtimmResource_i,
    rt_immMuxOutput_o
);


// Interface


// Calculate


endmodule
