module Control
(
    opCode_i,
    equal_i,
    branch_o,
    aluOP_o,
    aluSrc_o,
    memRead_o,
    memWrite_o,
    memToReg_o
);

// Interface

// Calculation

endmodule
