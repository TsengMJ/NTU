module Stall_MUX
(
    aluOp_i,
    aluSrc_i,
    memRead_i,
    memWrite_i,
    memToReg_i
    zero_i,

    aluOp_o,
    aluSrc_o,
    memRead_o,
    memWrite_o,
    memToReg_o
);

// Interface

// Calculate

endmodule
