module ALU_Input2_MUX
(
    rt_immMuxOutput_i,
    aluForwarding_i,
    memForwarding_i,
    forwardingB_i,
    aluInput2_o
);


// Interface


// Calculate


endmodule
