module
(
    aluOp_i,
    aluSrc_i,
    memRead_i,
    memWrite_i,
    memToReg_i,
    rsData_i,
    rtData_i,
    immExtended_i,
    rsAddr_i,
    rtAddr_i,
    rdAddr_i,

    aluOp_o,
    aluSrc_o,
    memRead_o,
    memWrite_o,
    memToReg_o,
    rsData_o,
    rtData_o,
    immExtended_o,
    rsAddr_o,
    rtAddr_o,
    rdAddr_o
);

// Interface

// Calculation


endmodule