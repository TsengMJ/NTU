module WB_MUX
(
    memData_i,
    aluResult_i,
    wbData_o
);

// Interface

// Calculate


endmodule
