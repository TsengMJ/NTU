module PC_Dst_MUX
(
    pcBranch_i,
    pcNext_i,
    pc_o
);

// Interface


// Calculate

endmodule
