module Register_MEM_WB
(
    memToReg_i,
    regWrite_i,
    memData_i,
    aluResult_i,
    wbAddr_i,

    memToReg_o,
    regWrite_o,
    memData_o,
    aluResult_o,
    wbAddr_o
);

// Interface

// Calculation

endmodule