module ALU_Input1_MUX
(
    rsData_i,
    aluForwarding_i,
    memForwarding_i,
    forwardingA_i,
    aluInput1_o
);


// Interface

// Calculate

endmodule
