module ALU
(
    aluInput1_i,
    aluInput2_i,
    aluCtrl_i,
    aluResult_o
);


// Interface


// Calculate


endmodule
