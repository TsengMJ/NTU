module Branch_Adder
(
    immShifted_i,
    instrAddr_i,
    pcBranch_o
);


// Interface


// Calculate


endmodule
