module Forwarding_Unit
(
    EX_rsAddr_i,
    EX_rtAddr_i,
    MEM_regWrite_i,
    MEM_wbAddr_i,
    WB_regWrite_i,
    WB_wbAddr_i,  

    forwardingA_o,
    forwardingB_o
);

// Interface

// Calculation

endmodule