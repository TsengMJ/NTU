module PC_Adder
(
    instrAddr_i,
    instrSize_i,
    pcNext_o
);

// Interface


// Calculation


endmodule
