module ALU_Ctrol
(
    funct_i,
    aluOp_i,
    aluCtrl_o

);

// Interface


// Calculate


endmodule
