module Shift
(
    immExtended_i,
    immShifted_o
);

// Interface


// Calculate


endmodule
