module Branch_Equal
(
    rsData_i,
    rtData_i,
    equal_o
);

// Interface


// Calculate


endmodule
